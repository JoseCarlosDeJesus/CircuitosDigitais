CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
30 140 1 210 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
12
13 Logic Switch~
5 388 362 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3536 0 0
2
5.89968e-315 0
0
6 74136~
219 215 431 0 3 22
0 5 4 2
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
4597 0 0
2
44212.5 0
0
6 74136~
219 215 385 0 3 22
0 6 4 3
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3835 0 0
2
44212.5 0
0
6 74136~
219 215 339 0 3 22
0 8 4 7
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3670 0 0
2
44212.5 0
0
6 74136~
219 218 282 0 3 22
0 10 4 9
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
5616 0 0
2
44212.5 0
0
14 Logic Display~
6 497 184 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 OF
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9323 0 0
2
5.89968e-315 0
0
14 Logic Display~
6 614 184 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 S1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
5.89968e-315 0
0
14 Logic Display~
6 591 184 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 S2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3108 0 0
2
5.89968e-315 0
0
14 Logic Display~
6 566 184 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 S3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4299 0 0
2
5.89968e-315 0
0
14 Logic Display~
6 543 184 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 S4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9672 0 0
2
5.89968e-315 0
0
6 74LS83
105 448 284 0 14 29
0 19 18 17 16 9 7 3 2 4
15 14 13 12 11
0
0 0 4848 0
6 74LS83
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
7876 0 0
2
5.89968e-315 0
0
9 Data Seq~
170 43 263 0 17 18
0 19 18 17 16 10 8 6 5 20
21 3 1 3 10 3 0 33
0
0 0 4720 0
6 DIGSRC
-21 -44 21 -36
3 DS1
-11 -44 10 -36
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
19 type:source { TW=1}
5 SIP10
21

0 8 7 6 5 4 3 2 1 9
10 8 7 6 5 4 3 2 1 9
10 0
65 0 0 512 1 0 0 0
2 DS
6369 0 0
2
5.89968e-315 0
0
AAJFABIJAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
22
3 8 2 0 0 4224 0 2 11 0 0 4
248 431
408 431
408 311
416 311
3 7 3 0 0 4224 0 3 11 0 0 4
248 385
408 385
408 302
416 302
0 2 4 0 0 8320 0 0 2 4 0 5
405 362
405 451
191 451
191 440
199 440
0 2 4 0 0 0 0 0 3 5 0 5
405 362
405 405
191 405
191 394
199 394
0 2 4 0 0 0 0 0 4 6 0 7
405 362
405 348
252 348
252 359
191 359
191 348
199 348
0 2 4 0 0 0 0 0 5 13 0 5
405 362
405 302
194 302
194 291
202 291
8 1 5 0 0 8320 0 12 2 0 0 4
75 299
181 299
181 422
199 422
7 1 6 0 0 4224 0 12 3 0 0 4
75 290
186 290
186 376
199 376
3 6 7 0 0 4224 0 4 11 0 0 4
248 339
403 339
403 293
416 293
6 1 8 0 0 4224 0 12 4 0 0 4
75 281
191 281
191 330
199 330
3 5 9 0 0 4224 0 5 11 0 0 4
251 282
408 282
408 284
416 284
5 1 10 0 0 4224 0 12 5 0 0 4
75 272
194 272
194 273
202 273
1 9 4 0 0 128 0 1 11 0 0 4
400 362
408 362
408 329
416 329
14 1 11 0 0 8320 0 11 6 0 0 3
481 329
497 329
497 202
13 1 12 0 0 4224 0 11 7 0 0 3
481 302
614 302
614 202
12 1 13 0 0 4224 0 11 8 0 0 3
481 293
591 293
591 202
11 1 14 0 0 4224 0 11 9 0 0 3
481 284
566 284
566 202
10 1 15 0 0 8320 0 11 10 0 0 3
481 275
543 275
543 202
4 4 16 0 0 4224 0 12 11 0 0 4
75 263
401 263
401 275
416 275
3 3 17 0 0 4224 0 12 11 0 0 4
75 254
401 254
401 266
416 266
2 2 18 0 0 4224 0 12 11 0 0 4
75 245
401 245
401 257
416 257
1 1 19 0 0 4224 0 12 11 0 0 4
75 236
401 236
401 248
416 248
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
