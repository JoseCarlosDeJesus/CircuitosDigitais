CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
10 0 30 50 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
18 D:\Circuit\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
70
13 Logic Switch~
5 187 1600 0 1 11
0 58
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 C
-2 -26 5 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
44273.9 10
0
13 Logic Switch~
5 197 1514 0 1 11
0 60
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 T0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
44273.9 9
0
13 Logic Switch~
5 195 1231 0 1 11
0 77
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 T7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
44273.9 8
0
13 Logic Switch~
5 196 1386 0 1 11
0 81
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 T3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
44273.9 7
0
13 Logic Switch~
5 196 1425 0 1 11
0 82
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 T2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
44273.9 6
0
13 Logic Switch~
5 197 1469 0 1 11
0 83
0
0 0 21360 0
2 0V
-4 -16 10 -8
2 T1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
44273.9 5
0
13 Logic Switch~
5 195 1349 0 1 11
0 80
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 T4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
44273.9 4
0
13 Logic Switch~
5 195 1312 0 1 11
0 79
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 T5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
44273.9 3
0
13 Logic Switch~
5 194 1275 0 1 11
0 78
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 T6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
44273.9 2
0
13 Logic Switch~
5 195 1193 0 1 11
0 76
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 T8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
44273.9 1
0
13 Logic Switch~
5 195 1153 0 1 11
0 75
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 T9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3472 0 0
2
44273.9 0
0
9 CA 7-Seg~
184 1320 1205 0 18 19
10 52 51 50 49 48 47 46 84 85
0 0 0 0 0 0 2 2 2
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
9998 0 0
2
44273.9 71
0
6 74LS47
187 1206 1456 0 14 29
0 8 10 12 14 86 87 46 47 48
49 50 51 52 88
0
0 0 4848 0
7 74LS247
-24 -60 25 -52
3 U19
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3536 0 0
2
44273.9 70
0
6 74LS47
187 1204 1678 0 14 29
0 7 9 11 13 89 90 39 40 41
42 43 44 45 91
0
0 0 4848 0
7 74LS247
-24 -60 25 -52
2 U5
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
4597 0 0
2
44273.9 69
0
12 D Flip-Flop~
219 925 1703 0 4 9
0 53 38 92 7
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U18
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3835 0 0
2
44273.9 68
0
12 D Flip-Flop~
219 925 1751 0 4 9
0 54 38 93 9
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U17
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3670 0 0
2
44273.9 67
0
12 D Flip-Flop~
219 926 1798 0 4 9
0 55 38 94 11
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U16
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
5616 0 0
2
44273.9 66
0
12 D Flip-Flop~
219 927 1846 0 4 9
0 56 38 95 13
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U15
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
9323 0 0
2
44273.9 65
0
12 D Flip-Flop~
219 928 1607 0 4 9
0 56 57 96 14
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U14
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
317 0 0
2
44273.9 64
0
12 D Flip-Flop~
219 927 1559 0 4 9
0 55 57 97 12
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U13
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3108 0 0
2
44273.9 63
0
12 D Flip-Flop~
219 926 1512 0 4 9
0 54 57 98 10
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U12
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
4299 0 0
2
44273.9 62
0
7 Ground~
168 783 1493 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9672 0 0
2
44273.9 61
0
5 4013~
219 714 1436 0 6 22
0 58 57 59 2 99 38
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U11B
19 -61 47 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 7 0
1 U
7876 0 0
2
44273.9 60
0
5 4013~
219 600 1436 0 6 22
0 2 38 59 58 100 57
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U11A
22 -61 50 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 3 0
1 U
6369 0 0
2
44273.9 59
0
12 D Flip-Flop~
219 926 1464 0 4 9
0 53 57 101 8
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U10
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
9172 0 0
2
44273.9 58
0
5 4071~
219 1026 1293 0 3 22
0 64 60 59
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U9A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
7100 0 0
2
44273.9 57
0
8 4-In OR~
219 931 1198 0 5 22
0 53 54 55 56 64
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U8A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 5 0
1 U
3820 0 0
2
44273.9 56
0
9 Inverter~
13 639 1249 0 2 22
0 61 56
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
7678 0 0
2
44273.9 55
0
9 Inverter~
13 639 1216 0 2 22
0 62 55
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
961 0 0
2
44273.9 54
0
9 Inverter~
13 638 1181 0 2 22
0 63 54
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
3178 0 0
2
44273.9 53
0
9 Inverter~
13 638 1148 0 2 22
0 65 53
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
3409 0 0
2
44273.9 52
0
5 74147
219 503 1166 0 13 27
0 66 67 68 69 70 71 72 73 74
61 62 63 65
0
0 0 4848 0
5 74147
-18 -60 17 -52
2 U6
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
121 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
27

0 10 5 4 3 2 1 13 12 11
9 7 6 14 10 5 4 3 2 1
13 12 11 9 7 6 14 0
65 0 0 0 1 0 0 0
1 U
3951 0 0
2
44273.9 51
0
9 Inverter~
13 267 1469 0 2 22
0 83 74
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
8885 0 0
2
44273.9 50
0
9 Inverter~
13 267 1425 0 2 22
0 82 73
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3780 0 0
2
44273.9 49
0
9 Inverter~
13 267 1386 0 2 22
0 81 72
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
9265 0 0
2
44273.9 48
0
9 Inverter~
13 267 1349 0 2 22
0 80 71
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
9442 0 0
2
44273.9 47
0
9 Inverter~
13 267 1312 0 2 22
0 79 70
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
9424 0 0
2
44273.9 46
0
9 Inverter~
13 267 1275 0 2 22
0 78 69
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
9968 0 0
2
44273.9 45
0
9 Inverter~
13 268 1231 0 2 22
0 77 68
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
9281 0 0
2
44273.9 44
0
9 Inverter~
13 267 1192 0 2 22
0 76 67
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
8464 0 0
2
44273.9 43
0
9 Inverter~
13 266 1153 0 2 22
0 75 66
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
7168 0 0
2
44273.9 42
0
9 CA 7-Seg~
184 1419 1205 0 18 19
10 45 44 43 42 41 40 39 102 103
0 0 0 0 0 0 2 2 2
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3171 0 0
2
44273.9 41
0
9 CA 7-Seg~
184 1827 1208 0 18 19
10 37 36 35 34 33 32 31 104 105
0 0 0 0 0 0 2 2 2
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP3
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
4139 0 0
2
44273.9 40
0
6 74LS47
187 1715 1453 0 14 29
0 3 4 5 6 106 107 31 32 33
34 35 36 37 108
0
0 0 4848 0
7 74LS247
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
6435 0 0
2
44273.9 37
0
7 Ground~
168 1263 203 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5283 0 0
2
44273.9 36
0
5 4071~
219 1533 237 0 3 22
0 29 28 24
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U9B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 6 0
1 U
6874 0 0
2
44273.9 35
0
5 4081~
219 1461 259 0 3 22
0 14 13 28
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U26B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 9 0
1 U
5305 0 0
2
44273.9 34
0
5 4081~
219 1461 215 0 3 22
0 30 2 29
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U26A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 9 0
1 U
34 0 0
2
44273.9 33
0
5 4030~
219 1403 163 0 3 22
0 30 2 6
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U25B
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 8 0
1 U
969 0 0
2
44273.9 32
0
5 4030~
219 1329 142 0 3 22
0 14 13 30
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U25A
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 8 0
1 U
8402 0 0
2
44273.9 31
0
5 4071~
219 1830 424 0 3 22
0 26 25 20
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U9D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 6 0
1 U
3751 0 0
2
44273.9 30
0
5 4081~
219 1758 446 0 3 22
0 12 11 25
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U27A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 10 0
1 U
4292 0 0
2
44273.9 29
0
5 4081~
219 1758 402 0 3 22
0 27 24 26
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U27B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 10 0
1 U
6118 0 0
2
44273.9 28
0
5 4030~
219 1700 350 0 3 22
0 27 24 5
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U28A
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 11 0
1 U
34 0 0
2
44273.9 27
0
5 4030~
219 1626 329 0 3 22
0 12 11 27
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U28B
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 11 0
1 U
6357 0 0
2
44273.9 26
0
5 4071~
219 2128 605 0 3 22
0 22 21 16
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U29A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 12 0
1 U
319 0 0
2
44273.9 25
0
5 4081~
219 2056 627 0 3 22
0 10 9 21
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U27C
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 10 0
1 U
3976 0 0
2
44273.9 24
0
5 4081~
219 2056 583 0 3 22
0 23 20 22
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U27D
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 10 0
1 U
7634 0 0
2
44273.9 23
0
5 4030~
219 1998 531 0 3 22
0 23 20 4
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U28C
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 11 0
1 U
523 0 0
2
44273.9 22
0
5 4030~
219 1924 510 0 3 22
0 10 9 23
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U28D
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 11 0
1 U
6748 0 0
2
44273.9 21
0
5 4071~
219 2451 800 0 3 22
0 18 17 15
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U29B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 12 0
1 U
6901 0 0
2
44273.9 20
0
5 4081~
219 2379 822 0 3 22
0 8 7 17
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U30A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 13 0
1 U
842 0 0
2
44273.9 19
0
5 4081~
219 2379 778 0 3 22
0 19 16 18
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U30B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 13 0
1 U
3277 0 0
2
44273.9 18
0
5 4030~
219 2321 726 0 3 22
0 19 16 3
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U31A
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 14 0
1 U
4212 0 0
2
44273.9 17
0
5 4030~
219 2247 705 0 3 22
0 8 7 19
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U31B
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 14 0
1 U
4720 0 0
2
44273.9 16
0
14 Logic Display~
6 2606 945 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5551 0 0
2
44273.9 15
0
14 Logic Display~
6 2634 946 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6986 0 0
2
44273.9 14
0
14 Logic Display~
6 2667 946 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8745 0 0
2
44273.9 13
0
14 Logic Display~
6 2703 944 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9592 0 0
2
44273.9 12
0
14 Logic Display~
6 2756 874 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8748 0 0
2
44273.9 11
0
138
1 0 3 0 0 12432 0 44 0 0 22 5
1683 1417
1674 1417
1674 1006
2619 1006
2619 963
2 0 4 0 0 12432 0 44 0 0 23 5
1683 1426
1670 1426
1670 1017
2650 1017
2650 961
3 0 5 0 0 12432 0 44 0 0 24 5
1683 1435
1663 1435
1663 1027
2689 1027
2689 964
4 0 6 0 0 12304 0 44 0 0 25 5
1683 1444
1659 1444
1659 1039
2712 1039
2712 962
0 2 7 0 0 8208 0 0 62 6 0 3
2173 714
2173 831
2355 831
2 0 7 0 0 4112 0 65 0 0 50 2
2231 714
1162 714
0 1 8 0 0 8208 0 0 62 8 0 3
2188 696
2188 813
2355 813
1 0 8 0 0 4112 0 65 0 0 54 2
2231 696
1119 696
2 0 9 0 0 4112 0 57 0 0 10 3
2032 636
1844 636
1844 519
2 0 9 0 0 4112 0 60 0 0 51 2
1908 519
1153 519
1 0 10 0 0 4112 0 57 0 0 12 3
2032 618
1855 618
1855 501
1 0 10 0 0 4112 0 60 0 0 55 2
1908 501
1108 501
0 2 11 0 0 8208 0 0 52 14 0 3
1564 338
1564 455
1734 455
2 0 11 0 0 4112 0 55 0 0 52 2
1610 338
1145 338
0 1 12 0 0 8208 0 0 52 16 0 3
1576 320
1576 437
1734 437
1 0 12 0 0 4112 0 55 0 0 56 2
1610 320
1097 320
0 2 13 0 0 8208 0 0 47 18 0 3
1284 151
1284 268
1437 268
2 0 13 0 0 4112 0 50 0 0 53 2
1313 151
1136 151
1 0 14 0 0 4112 0 47 0 0 20 3
1437 250
1295 250
1295 133
1 0 14 0 0 4112 0 50 0 0 57 2
1313 133
1086 133
3 1 15 0 0 8336 0 61 70 0 0 3
2484 800
2484 892
2756 892
1 3 3 0 0 16 0 66 64 0 0 4
2606 963
2620 963
2620 726
2354 726
3 1 4 0 0 16 0 59 67 0 0 4
2031 531
2650 531
2650 964
2634 964
1 3 5 0 0 16 0 68 54 0 0 4
2667 964
2689 964
2689 350
1733 350
3 1 6 0 0 4240 0 49 69 0 0 4
1436 163
2712 163
2712 962
2703 962
0 2 16 0 0 8336 0 0 63 27 0 3
2201 735
2201 787
2355 787
3 2 16 0 0 16 0 56 64 0 0 4
2161 605
2201 605
2201 735
2305 735
3 2 17 0 0 12432 0 62 61 0 0 4
2400 822
2414 822
2414 809
2438 809
3 1 18 0 0 12432 0 63 61 0 0 4
2400 778
2414 778
2414 791
2438 791
0 1 19 0 0 8336 0 0 63 31 0 3
2294 717
2294 769
2355 769
3 1 19 0 0 16 0 65 64 0 0 4
2280 705
2294 705
2294 717
2305 717
0 2 20 0 0 8336 0 0 58 33 0 3
1871 540
1871 592
2032 592
3 2 20 0 0 16 0 51 59 0 0 4
1863 424
1871 424
1871 540
1982 540
3 2 21 0 0 12432 0 57 56 0 0 4
2077 627
2091 627
2091 614
2115 614
3 1 22 0 0 12432 0 58 56 0 0 4
2077 583
2091 583
2091 596
2115 596
0 1 23 0 0 8336 0 0 58 37 0 3
1971 522
1971 574
2032 574
3 1 23 0 0 16 0 60 59 0 0 4
1957 510
1971 510
1971 522
1982 522
0 2 24 0 0 8336 0 0 53 39 0 3
1588 359
1588 411
1734 411
3 2 24 0 0 16 0 46 54 0 0 4
1566 237
1588 237
1588 359
1684 359
3 2 25 0 0 12432 0 52 51 0 0 4
1779 446
1793 446
1793 433
1817 433
3 1 26 0 0 12432 0 53 51 0 0 4
1779 402
1793 402
1793 415
1817 415
0 1 27 0 0 8336 0 0 53 43 0 3
1673 341
1673 393
1734 393
3 1 27 0 0 16 0 55 54 0 0 4
1659 329
1673 329
1673 341
1684 341
3 2 28 0 0 12432 0 47 46 0 0 4
1482 259
1496 259
1496 246
1520 246
3 1 29 0 0 12432 0 48 46 0 0 4
1482 215
1496 215
1496 228
1520 228
0 2 2 0 0 8208 0 0 48 47 0 3
1338 172
1338 224
1437 224
2 1 2 0 0 4112 0 49 45 0 0 3
1387 172
1263 172
1263 197
0 1 30 0 0 8336 0 0 48 49 0 3
1376 154
1376 206
1437 206
3 1 30 0 0 16 0 50 49 0 0 4
1362 142
1376 142
1376 154
1387 154
0 0 7 0 0 4240 0 0 0 0 83 4
1162 105
1162 1627
1160 1627
1160 1642
0 0 9 0 0 4240 0 0 0 0 80 4
1153 106
1153 1636
1151 1636
1151 1651
0 0 11 0 0 4240 0 0 0 0 81 4
1145 106
1145 1645
1141 1645
1141 1660
0 0 13 0 0 4240 0 0 0 0 82 4
1136 105
1136 1654
1131 1654
1131 1669
0 0 8 0 0 4240 0 0 0 87 0 2
1119 1420
1119 109
0 0 10 0 0 4240 0 0 0 84 0 4
1108 1429
1108 350
1107 350
1107 110
0 0 12 0 0 4240 0 0 0 85 0 4
1098 1438
1098 359
1097 359
1097 112
0 0 14 0 0 4240 0 0 0 86 0 2
1086 1447
1086 113
7 7 31 0 0 8336 0 44 43 0 0 3
1753 1417
1842 1417
1842 1244
8 6 32 0 0 8336 0 44 43 0 0 3
1753 1426
1836 1426
1836 1244
9 5 33 0 0 8336 0 44 43 0 0 3
1753 1435
1830 1435
1830 1244
10 4 34 0 0 8336 0 44 43 0 0 3
1753 1444
1824 1444
1824 1244
11 3 35 0 0 8336 0 44 43 0 0 3
1753 1453
1818 1453
1818 1244
12 2 36 0 0 8336 0 44 43 0 0 3
1753 1462
1812 1462
1812 1244
13 1 37 0 0 8336 0 44 43 0 0 3
1753 1471
1806 1471
1806 1244
6 0 38 0 0 4112 0 23 0 0 103 2
738 1400
807 1400
7 7 39 0 0 4240 0 42 14 0 0 3
1434 1241
1434 1642
1242 1642
6 8 40 0 0 4240 0 42 14 0 0 3
1428 1241
1428 1651
1242 1651
5 9 41 0 0 4240 0 42 14 0 0 3
1422 1241
1422 1660
1242 1660
4 10 42 0 0 4240 0 42 14 0 0 3
1416 1241
1416 1669
1242 1669
3 11 43 0 0 4240 0 42 14 0 0 3
1410 1241
1410 1678
1242 1678
2 12 44 0 0 4240 0 42 14 0 0 3
1404 1241
1404 1687
1242 1687
1 13 45 0 0 4240 0 42 14 0 0 3
1398 1241
1398 1696
1242 1696
7 7 46 0 0 4240 0 12 13 0 0 3
1335 1241
1335 1420
1244 1420
6 8 47 0 0 4240 0 12 13 0 0 3
1329 1241
1329 1429
1244 1429
5 9 48 0 0 4240 0 12 13 0 0 3
1323 1241
1323 1438
1244 1438
4 10 49 0 0 4240 0 12 13 0 0 3
1317 1241
1317 1447
1244 1447
3 11 50 0 0 4240 0 12 13 0 0 3
1311 1241
1311 1456
1244 1456
2 12 51 0 0 4240 0 12 13 0 0 3
1305 1241
1305 1465
1244 1465
1 13 52 0 0 4240 0 12 13 0 0 3
1299 1241
1299 1474
1244 1474
4 2 9 0 0 16 0 16 14 0 0 4
949 1715
1038 1715
1038 1651
1172 1651
4 3 11 0 0 16 0 17 14 0 0 4
950 1762
1047 1762
1047 1660
1172 1660
4 4 13 0 0 16 0 18 14 0 0 4
951 1810
1056 1810
1056 1669
1172 1669
4 1 7 0 0 16 0 15 14 0 0 4
949 1667
964 1667
964 1642
1172 1642
4 2 10 0 0 16 0 21 13 0 0 4
950 1476
1020 1476
1020 1429
1174 1429
4 3 12 0 0 16 0 20 13 0 0 4
951 1523
1032 1523
1032 1438
1174 1438
4 4 14 0 0 16 0 19 13 0 0 4
952 1571
1047 1571
1047 1447
1174 1447
4 1 8 0 0 16 0 25 13 0 0 4
950 1428
965 1428
965 1420
1174 1420
1 0 53 0 0 4112 0 25 0 0 92 2
902 1428
890 1428
1 0 54 0 0 4112 0 21 0 0 93 2
902 1476
876 1476
1 0 55 0 0 4112 0 20 0 0 94 2
903 1523
860 1523
1 0 56 0 0 4112 0 19 0 0 95 2
904 1571
845 1571
1 0 53 0 0 8336 0 15 0 0 116 3
901 1667
890 1667
890 1185
1 0 54 0 0 8336 0 16 0 0 118 3
901 1715
876 1715
876 1194
1 0 55 0 0 8336 0 17 0 0 119 3
902 1762
860 1762
860 1203
1 0 56 0 0 8336 0 18 0 0 117 3
903 1810
845 1810
845 1212
2 0 57 0 0 4112 0 20 0 0 98 2
903 1541
831 1541
2 0 57 0 0 16 0 21 0 0 98 2
902 1494
831 1494
2 0 57 0 0 8208 0 25 0 0 99 3
902 1446
831 1446
831 1589
0 2 57 0 0 8336 0 0 19 106 0 3
649 1400
649 1589
904 1589
2 0 38 0 0 4112 0 15 0 0 103 2
901 1685
807 1685
2 0 38 0 0 16 0 16 0 0 103 2
901 1733
807 1733
2 0 38 0 0 4112 0 17 0 0 103 2
902 1780
807 1780
2 2 38 0 0 16528 0 24 18 0 0 6
576 1400
564 1400
564 1350
807 1350
807 1828
903 1828
4 0 58 0 0 4112 0 24 0 0 105 2
600 1442
600 1600
1 1 58 0 0 16528 0 23 1 0 0 5
714 1379
714 1372
682 1372
682 1600
199 1600
6 2 57 0 0 16 0 24 23 0 0 2
624 1400
690 1400
4 0 2 0 0 16 0 23 0 0 108 3
714 1442
714 1469
783 1469
1 1 2 0 0 8336 0 24 22 0 0 4
600 1379
600 1362
783 1362
783 1487
3 0 59 0 0 8208 0 23 0 0 110 3
690 1418
671 1418
671 1334
3 3 59 0 0 12432 0 26 24 0 0 6
1059 1293
1079 1293
1079 1334
527 1334
527 1418
576 1418
2 1 60 0 0 4240 0 26 2 0 0 4
1013 1302
477 1302
477 1514
209 1514
10 1 61 0 0 8336 0 32 28 0 0 4
541 1175
599 1175
599 1249
624 1249
11 1 62 0 0 4240 0 32 29 0 0 4
541 1166
608 1166
608 1216
624 1216
12 1 63 0 0 4240 0 32 30 0 0 4
541 1157
616 1157
616 1181
623 1181
5 1 64 0 0 8336 0 27 26 0 0 4
964 1198
991 1198
991 1284
1013 1284
2 1 53 0 0 16 0 31 27 0 0 4
659 1148
684 1148
684 1185
914 1185
2 4 56 0 0 16 0 28 27 0 0 4
660 1249
684 1249
684 1212
914 1212
2 2 54 0 0 16 0 30 27 0 0 4
659 1181
677 1181
677 1194
914 1194
2 3 55 0 0 16 0 29 27 0 0 4
660 1216
677 1216
677 1203
914 1203
13 1 65 0 0 4240 0 32 31 0 0 2
541 1148
623 1148
2 1 66 0 0 4240 0 41 32 0 0 4
287 1153
378 1153
378 1130
465 1130
2 2 67 0 0 4240 0 40 32 0 0 4
288 1192
388 1192
388 1139
465 1139
2 3 68 0 0 4240 0 39 32 0 0 4
289 1231
399 1231
399 1148
465 1148
2 4 69 0 0 4240 0 38 32 0 0 4
288 1275
409 1275
409 1157
465 1157
2 5 70 0 0 8336 0 37 32 0 0 4
288 1312
419 1312
419 1166
465 1166
2 6 71 0 0 8336 0 36 32 0 0 4
288 1349
430 1349
430 1175
465 1175
2 7 72 0 0 8336 0 35 32 0 0 4
288 1386
443 1386
443 1184
465 1184
2 8 73 0 0 8336 0 34 32 0 0 4
288 1425
455 1425
455 1193
465 1193
2 9 74 0 0 8336 0 33 32 0 0 3
288 1469
465 1469
465 1202
1 1 75 0 0 4240 0 11 41 0 0 2
207 1153
251 1153
1 1 76 0 0 8336 0 10 40 0 0 3
207 1193
207 1192
252 1192
1 1 77 0 0 4240 0 3 39 0 0 2
207 1231
253 1231
1 1 78 0 0 4240 0 9 38 0 0 2
206 1275
252 1275
1 1 79 0 0 4240 0 8 37 0 0 2
207 1312
252 1312
1 1 80 0 0 4240 0 7 36 0 0 2
207 1349
252 1349
1 1 81 0 0 4240 0 4 35 0 0 2
208 1386
252 1386
1 1 82 0 0 4240 0 5 34 0 0 2
208 1425
252 1425
1 1 83 0 0 4240 0 6 33 0 0 2
209 1469
252 1469
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
