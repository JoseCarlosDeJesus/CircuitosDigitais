CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
20 110 30 150 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
27
13 Logic Switch~
5 193 681 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3215 0 0
2
44183.6 0
0
13 Logic Switch~
5 195 616 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7903 0 0
2
44183.6 0
0
13 Logic Switch~
5 195 563 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7121 0 0
2
44183.6 0
0
13 Logic Switch~
5 198 509 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4484 0 0
2
44183.6 0
0
13 Logic Switch~
5 279 347 0 1 11
0 20
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5996 0 0
2
5.89966e-315 0
0
13 Logic Switch~
5 313 234 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7804 0 0
2
5.89966e-315 0
0
13 Logic Switch~
5 315 183 0 1 11
0 21
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5523 0 0
2
5.89966e-315 0
0
13 Logic Switch~
5 319 134 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3330 0 0
2
5.89966e-315 0
0
14 Logic Display~
6 651 503 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3465 0 0
2
44183.6 0
0
8 2-In OR~
219 550 580 0 3 22
0 3 4 2
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
8396 0 0
2
44183.6 0
0
5 7415~
219 437 575 0 4 22
0 7 5 6 3
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 7 0
1 U
3685 0 0
2
44183.6 0
0
9 Inverter~
13 282 677 0 2 22
0 8 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 6 0
1 U
7849 0 0
2
44183.6 0
0
9 Inverter~
13 282 509 0 2 22
0 9 7
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 6 0
1 U
6343 0 0
2
44183.6 0
0
9 Inverter~
13 260 563 0 2 22
0 5 11
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
7376 0 0
2
44183.6 0
0
9 2-In AND~
219 333 577 0 3 22
0 11 10 4
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
9156 0 0
2
44183.6 0
0
14 Logic Display~
6 758 213 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5776 0 0
2
5.89966e-315 0
0
8 3-In OR~
219 623 275 0 4 22
0 13 14 15 12
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U4A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 4 0
1 U
7207 0 0
2
5.89966e-315 0
0
9 Inverter~
13 409 410 0 2 22
0 18 19
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
4459 0 0
2
5.89966e-315 0
0
5 7415~
219 453 419 0 4 22
0 19 16 17 15
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 1 0
1 U
3760 0 0
2
5.89966e-315 0
0
9 Inverter~
13 367 418 0 2 22
0 22 17
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
754 0 0
2
5.89966e-315 0
0
9 Inverter~
13 293 408 0 2 22
0 18 23
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
9767 0 0
2
5.89966e-315 0
0
5 7415~
219 336 417 0 4 22
0 23 21 20 22
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 1 0
1 U
7978 0 0
2
5.89966e-315 0
0
9 Inverter~
13 397 304 0 2 22
0 18 24
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
3142 0 0
2
5.89966e-315 0
0
9 Inverter~
13 369 322 0 2 22
0 16 25
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
3284 0 0
2
5.89966e-315 0
0
9 4-In AND~
219 457 317 0 5 22
0 24 21 25 20 14
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U3A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 3 0
1 U
659 0 0
2
5.89966e-315 0
0
9 Inverter~
13 371 183 0 2 22
0 21 26
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
3800 0 0
2
5.89966e-315 0
0
5 7415~
219 453 195 0 4 22
0 18 26 16 13
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 1 0
1 U
6792 0 0
2
5.89966e-315 0
0
34
3 1 2 0 0 4224 0 10 9 0 0 3
583 580
651 580
651 521
4 1 3 0 0 4224 0 11 10 0 0 4
458 575
529 575
529 571
537 571
3 2 4 0 0 12416 0 15 10 0 0 6
354 577
409 577
409 595
529 595
529 589
537 589
0 2 5 0 0 8320 0 0 11 11 0 5
225 563
225 597
400 597
400 575
413 575
2 3 6 0 0 4224 0 12 11 0 0 4
303 677
405 677
405 584
413 584
2 1 7 0 0 4224 0 13 11 0 0 4
303 509
405 509
405 566
413 566
1 1 8 0 0 4224 0 1 12 0 0 4
205 681
259 681
259 677
267 677
1 1 9 0 0 4224 0 4 13 0 0 2
210 509
267 509
1 2 10 0 0 4224 0 2 15 0 0 4
207 616
301 616
301 586
309 586
2 1 11 0 0 4224 0 14 15 0 0 4
281 563
301 563
301 568
309 568
1 1 5 0 0 0 0 3 14 0 0 2
207 563
245 563
4 1 12 0 0 4224 0 17 16 0 0 3
656 275
758 275
758 231
4 1 13 0 0 4224 0 27 17 0 0 4
474 195
602 195
602 266
610 266
5 2 14 0 0 4224 0 25 17 0 0 4
478 317
597 317
597 275
611 275
4 3 15 0 0 8320 0 19 17 0 0 4
474 419
602 419
602 284
610 284
0 2 16 0 0 4224 0 0 19 32 0 3
395 234
395 419
429 419
2 3 17 0 0 8320 0 20 19 0 0 3
388 418
388 428
429 428
0 1 18 0 0 4224 0 0 18 34 0 3
373 134
373 410
394 410
2 1 19 0 0 4224 0 18 19 0 0 2
430 410
429 410
0 3 20 0 0 4096 0 0 22 25 0 3
304 347
304 426
312 426
1 2 21 0 0 4224 0 7 22 0 0 3
327 183
327 417
312 417
0 1 18 0 0 0 0 0 21 34 0 5
336 134
336 393
270 393
270 408
278 408
1 4 22 0 0 8320 0 20 22 0 0 3
352 418
352 417
357 417
2 1 23 0 0 4224 0 21 22 0 0 2
314 408
312 408
1 4 20 0 0 4224 0 5 25 0 0 4
291 347
425 347
425 331
433 331
2 1 24 0 0 4224 0 23 25 0 0 2
418 304
433 304
2 3 25 0 0 4224 0 24 25 0 0 2
390 322
433 322
0 1 16 0 0 0 0 0 24 32 0 3
334 234
334 322
354 322
0 2 21 0 0 0 0 0 25 33 0 3
341 183
341 313
433 313
0 1 18 0 0 0 0 0 23 34 0 3
351 134
351 304
382 304
2 2 26 0 0 4224 0 26 27 0 0 4
392 183
416 183
416 195
429 195
1 3 16 0 0 0 0 6 27 0 0 4
325 234
421 234
421 204
429 204
1 1 21 0 0 0 0 7 26 0 0 2
327 183
356 183
1 1 18 0 0 0 0 8 27 0 0 4
331 134
421 134
421 186
429 186
10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
306 451 457 475
313 457 449 473
17 Circuito Reduzido
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
229 649 252 673
236 655 244 671
1 D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
225 591 248 615
232 596 240 612
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
221 533 244 557
228 538 236 554
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
218 461 241 485
225 467 233 483
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
331 153 354 177
338 158 346 174
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
340 109 363 133
347 115 355 131
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
336 211 359 235
343 217 351 233
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
303 323 326 347
310 328 318 344
1 D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
380 77 563 101
387 82 555 98
21 Circuito N�o Reduzido
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
