CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 460 1 110 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
27
13 Logic Switch~
5 1235 1154 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7678 0 0
2
5.89975e-315 0
0
8 2-In OR~
219 779 752 0 3 22
0 10 9 11
0
0 0 624 512
6 74LS32
-21 -24 21 -16
4 U12A
-2 -25 26 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
961 0 0
2
5.89975e-315 5.26354e-315
0
8 3-In OR~
219 744 574 0 4 22
0 6 7 8 12
0
0 0 624 512
4 4075
-14 -24 14 -16
4 U14A
-2 -25 26 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 10 0
1 U
3178 0 0
2
5.89975e-315 5.30499e-315
0
5 7415~
219 916 795 0 4 22
0 5 5 5 9
0
0 0 624 512
6 74LS15
-21 -28 21 -20
4 U13B
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 9 0
1 U
3409 0 0
2
5.89975e-315 5.32571e-315
0
5 7415~
219 920 757 0 4 22
0 5 5 5 10
0
0 0 624 512
6 74LS15
-21 -28 21 -20
4 U13A
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 9 0
1 U
3951 0 0
2
5.89975e-315 5.34643e-315
0
9 2-In AND~
219 919 680 0 3 22
0 5 5 8
0
0 0 624 512
6 74LS08
-21 -24 21 -16
4 U11A
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
8885 0 0
2
5.89975e-315 5.3568e-315
0
9 2-In AND~
219 914 632 0 3 22
0 5 5 7
0
0 0 624 512
6 74LS08
-21 -24 21 -16
3 U9D
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3780 0 0
2
5.89975e-315 5.36716e-315
0
9 2-In AND~
219 911 572 0 3 22
0 5 5 6
0
0 0 624 512
6 74LS08
-21 -24 21 -16
3 U9C
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
9265 0 0
2
5.89975e-315 5.37752e-315
0
9 Inverter~
13 625 801 0 2 22
0 11 13
0
0 0 624 512
6 74LS04
-21 -19 21 -11
3 U7C
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
9442 0 0
2
5.89975e-315 5.38788e-315
0
9 2-In NOR~
219 484 924 0 3 22
0 12 11 2
0
0 0 624 180
6 74LS02
-21 -24 21 -16
4 U10A
4 -25 32 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
9424 0 0
2
5.89975e-315 5.39306e-315
0
9 2-In AND~
219 483 810 0 3 22
0 12 13 4
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U9B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
9968 0 0
2
5.89975e-315 5.39824e-315
0
9 2-In AND~
219 443 741 0 3 22
0 12 11 3
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U9A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
9281 0 0
2
5.89975e-315 5.40342e-315
0
9 Inverter~
13 525 1016 0 2 22
0 4 14
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
8464 0 0
2
5.89975e-315 5.4086e-315
0
7 Buffer~
58 412 1063 0 2 22
0 2 15
0
0 0 624 0
4 4050
-14 -19 14 -11
3 U6B
-11 -20 10 -12
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
7168 0 0
2
5.89975e-315 5.41378e-315
0
6 74266~
219 659 1044 0 3 22
0 3 15 16
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U8A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3171 0 0
2
5.89975e-315 5.41896e-315
0
9 Inverter~
13 1154 908 0 2 22
0 22 5
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U7A
12 -18 33 -10
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
4139 0 0
2
5.89975e-315 5.42414e-315
0
7 Buffer~
58 1120 878 0 2 22
0 22 5
0
0 0 624 90
4 4050
-14 -19 14 -11
3 U6A
2 -22 23 -14
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
6435 0 0
2
5.89975e-315 5.42933e-315
0
7 Buffer~
58 1091 836 0 2 22
0 21 5
0
0 0 624 90
4 4050
-14 -19 14 -11
3 U5F
4 -20 25 -12
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
5283 0 0
2
5.89975e-315 5.43192e-315
0
7 Buffer~
58 1062 916 0 2 22
0 20 5
0
0 0 624 90
4 4050
-14 -19 14 -11
3 U5D
8 -17 29 -9
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
6874 0 0
2
5.89975e-315 5.43451e-315
0
7 Buffer~
58 1030 884 0 2 22
0 19 5
0
0 0 624 90
4 4050
-14 -19 14 -11
3 U5C
1 -18 22 -10
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
5305 0 0
2
5.89975e-315 5.4371e-315
0
7 Buffer~
58 993 862 0 2 22
0 23 5
0
0 0 624 90
4 4050
-14 -19 14 -11
3 U5A
4 -21 25 -13
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
34 0 0
2
5.89975e-315 5.43969e-315
0
12 D Flip-Flop~
219 902 896 0 4 9
0 12 18 24 20
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U4
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
969 0 0
2
5.89975e-315 5.44228e-315
0
12 D Flip-Flop~
219 900 951 0 4 9
0 11 18 19 23
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U3
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
8402 0 0
2
5.89975e-315 5.44487e-315
0
4 4024
219 921 1011 0 9 19
0 17 16 25 26 27 22 28 29 30
0
0 0 4848 0
4 4024
-14 -60 14 -52
2 U2
-7 -61 7 -53
0
15 DVDD=14;DGND=7;
69 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 1 2 12 11 9 6 5 4 3
1 2 12 11 9 6 5 4 3 0
65 0 0 512 1 0 0 0
1 U
3751 0 0
2
5.89975e-315 5.44746e-315
0
4 4024
219 1038 1067 0 9 19
0 17 14 31 32 21 33 34 35 36
0
0 0 4848 0
4 4024
-14 -60 14 -52
2 U1
-7 -61 7 -53
0
15 DVDD=14;DGND=7;
69 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 1 2 12 11 9 6 5 4 3
1 2 12 11 9 6 5 4 3 0
65 0 0 512 1 0 0 0
1 U
4292 0 0
2
5.89975e-315 5.45005e-315
0
10 StopLight~
181 209 1143 0 10 13
0 3 4 2 0 0 0 0 0 0
1
0
0 0 21088 512
4 1MEG
-15 -42 13 -34
4 SEM1
-20 -34 8 -26
0
0
37 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
0
0
0
7

0 1 2 3 1 2 3 0
82 0 0 0 1 0 0 0
3 SEM
6118 0 0
2
5.89975e-315 5.45264e-315
0
7 Pulser~
4 626 1222 0 10 12
0 37 38 17 18 0 0 50 50 44
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 1 0 0
1 V
34 0 0
2
5.89975e-315 5.45523e-315
0
51
1 0 2 0 0 4224 0 14 0 0 4 3
397 1063
330 1063
330 1019
1 0 3 0 0 4224 0 15 0 0 6 3
643 1035
383 1035
383 864
1 0 4 0 0 8320 0 13 0 0 5 3
510 1016
453 1016
453 932
3 3 2 0 0 16512 0 10 26 0 0 5
457 924
330 924
330 1019
219 1019
219 1157
3 2 4 0 0 16512 0 11 26 0 0 6
456 810
453 810
453 932
295 932
295 1143
219 1143
3 1 3 0 0 16512 0 12 26 0 0 6
416 741
383 741
383 864
260 864
260 1129
219 1129
3 0 5 0 0 4096 0 4 0 0 51 2
936 804
997 804
2 0 5 0 0 4096 0 4 0 0 48 4
936 795
1041 795
1041 794
1056 794
1 0 5 0 0 4096 0 4 0 0 45 4
936 786
1140 786
1140 785
1155 785
1 0 5 0 0 0 0 5 0 0 47 4
940 748
1086 748
1086 708
1101 708
2 0 5 0 0 0 0 5 0 0 48 4
940 757
1041 757
1041 717
1056 717
3 0 5 0 0 0 0 5 0 0 49 4
940 766
1013 766
1013 726
1028 726
2 0 5 0 0 0 0 6 0 0 49 4
939 689
1013 689
1013 655
1028 655
1 0 5 0 0 4096 0 6 0 0 51 4
939 671
1250 671
1250 637
1420 637
2 0 5 0 0 0 0 7 0 0 49 4
934 641
1008 641
1008 595
1028 595
1 0 5 0 0 0 0 7 0 0 46 4
934 623
1117 623
1117 578
1132 578
2 0 5 0 0 0 0 8 0 0 48 4
931 581
1041 581
1041 529
1056 529
1 0 5 0 0 0 0 8 0 0 45 4
931 563
1140 563
1140 511
1155 511
1 3 6 0 0 4224 0 3 8 0 0 4
763 565
840 565
840 572
886 572
2 3 7 0 0 4224 0 3 7 0 0 4
762 574
851 574
851 632
889 632
3 3 8 0 0 8320 0 3 6 0 0 4
763 583
859 583
859 680
894 680
2 4 9 0 0 12416 0 2 4 0 0 4
798 761
838 761
838 795
891 795
1 4 10 0 0 4224 0 2 5 0 0 4
798 743
855 743
855 757
895 757
2 0 11 0 0 4096 0 10 0 0 30 3
509 915
741 915
741 873
1 0 11 0 0 0 0 9 0 0 30 4
646 801
726 801
726 859
741 859
2 0 11 0 0 4224 0 12 0 0 30 4
461 732
726 732
726 800
741 800
1 0 12 0 0 4096 0 12 0 0 31 4
461 750
687 750
687 818
702 818
1 0 12 0 0 0 0 11 0 0 31 4
501 819
670 819
670 877
702 877
1 0 12 0 0 0 0 10 0 0 31 4
509 933
679 933
679 932
702 932
1 3 11 0 0 128 0 23 2 0 0 5
876 915
741 915
741 800
752 800
752 752
1 4 12 0 0 16512 0 22 3 0 0 6
878 860
702 860
702 932
702 932
702 574
717 574
2 2 13 0 0 4224 0 11 9 0 0 2
501 801
610 801
2 2 14 0 0 4224 0 25 13 0 0 4
1006 1076
563 1076
563 1016
546 1016
2 2 15 0 0 12416 0 15 14 0 0 4
643 1053
566 1053
566 1063
427 1063
2 3 16 0 0 12416 0 24 15 0 0 4
889 1020
879 1020
879 1044
698 1044
0 1 17 0 0 12288 0 0 24 37 0 4
816 1120
816 1177
883 1177
883 1002
3 1 17 0 0 8336 0 27 25 0 0 9
650 1213
650 1217
1002 1217
1002 1151
912 1151
912 1131
816 1131
816 1058
1000 1058
0 2 18 0 0 4096 0 0 22 39 0 3
840 952
840 878
878 878
4 2 18 0 0 8320 0 27 23 0 0 9
656 1222
656 1220
996 1220
996 1160
906 1160
906 1140
840 1140
840 933
876 933
1 3 19 0 0 8320 0 20 23 0 0 3
1030 899
1030 933
930 933
1 4 20 0 0 8320 0 19 22 0 0 3
1062 931
1062 860
926 860
1 5 21 0 0 4224 0 18 25 0 0 3
1091 851
1091 1067
1070 1067
1 0 22 0 0 4096 0 16 0 0 44 3
1157 926
1157 1020
1132 1020
1 6 22 0 0 16512 0 17 24 0 0 5
1120 893
1120 1020
1132 1020
1132 1002
953 1002
0 2 5 0 0 0 0 0 16 51 0 4
1155 511
1155 785
1157 785
1157 890
0 2 5 0 0 0 0 0 17 51 0 4
1132 511
1132 578
1120 578
1120 863
0 2 5 0 0 0 0 0 18 51 0 4
1101 511
1101 708
1091 708
1091 821
0 2 5 0 0 0 0 0 19 51 0 4
1056 511
1056 794
1062 794
1062 901
0 2 5 0 0 0 0 0 20 51 0 4
1028 511
1028 726
1030 726
1030 869
1 4 23 0 0 8320 0 21 23 0 0 3
993 877
993 915
924 915
1 2 5 0 0 8320 0 1 21 0 0 7
1247 1154
1420 1154
1420 511
997 511
997 804
993 804
993 847
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
